module memory_game();

endmodule
